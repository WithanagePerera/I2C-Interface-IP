// IMPORTANT: This is the address of the I2C slave
localparam I2C_ADDR = 7'b0001000;
